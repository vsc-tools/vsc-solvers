
package vsc_solvers;
    `include "vsc_constraint_set.svh"

    `include "vsc_expr.svh"
    `include "vsc_expr_bit.svh"
    `include "vsc_expr_lt_u.svh"
    `include "vsc_expr_zext.svh"

    `include "vsc_if_else.svh"


endpackage

