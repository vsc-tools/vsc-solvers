
class VscVarBit;
endclass
